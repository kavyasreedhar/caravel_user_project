magic
tech sky130A
magscale 1 2
timestamp 1622790553
<< obsli1 >>
rect 1104 1377 178848 117521
<< obsm1 >>
rect 106 348 179846 117552
<< metal2 >>
rect 754 119200 810 120000
rect 2318 119200 2374 120000
rect 3882 119200 3938 120000
rect 5446 119200 5502 120000
rect 7010 119200 7066 120000
rect 8574 119200 8630 120000
rect 10230 119200 10286 120000
rect 11794 119200 11850 120000
rect 13358 119200 13414 120000
rect 14922 119200 14978 120000
rect 16486 119200 16542 120000
rect 18050 119200 18106 120000
rect 19706 119200 19762 120000
rect 21270 119200 21326 120000
rect 22834 119200 22890 120000
rect 24398 119200 24454 120000
rect 25962 119200 26018 120000
rect 27526 119200 27582 120000
rect 29182 119200 29238 120000
rect 30746 119200 30802 120000
rect 32310 119200 32366 120000
rect 33874 119200 33930 120000
rect 35438 119200 35494 120000
rect 37002 119200 37058 120000
rect 38658 119200 38714 120000
rect 40222 119200 40278 120000
rect 41786 119200 41842 120000
rect 43350 119200 43406 120000
rect 44914 119200 44970 120000
rect 46478 119200 46534 120000
rect 48134 119200 48190 120000
rect 49698 119200 49754 120000
rect 51262 119200 51318 120000
rect 52826 119200 52882 120000
rect 54390 119200 54446 120000
rect 55954 119200 56010 120000
rect 57610 119200 57666 120000
rect 59174 119200 59230 120000
rect 60738 119200 60794 120000
rect 62302 119200 62358 120000
rect 63866 119200 63922 120000
rect 65430 119200 65486 120000
rect 67086 119200 67142 120000
rect 68650 119200 68706 120000
rect 70214 119200 70270 120000
rect 71778 119200 71834 120000
rect 73342 119200 73398 120000
rect 74906 119200 74962 120000
rect 76562 119200 76618 120000
rect 78126 119200 78182 120000
rect 79690 119200 79746 120000
rect 81254 119200 81310 120000
rect 82818 119200 82874 120000
rect 84382 119200 84438 120000
rect 86038 119200 86094 120000
rect 87602 119200 87658 120000
rect 89166 119200 89222 120000
rect 90730 119200 90786 120000
rect 92294 119200 92350 120000
rect 93858 119200 93914 120000
rect 95514 119200 95570 120000
rect 97078 119200 97134 120000
rect 98642 119200 98698 120000
rect 100206 119200 100262 120000
rect 101770 119200 101826 120000
rect 103334 119200 103390 120000
rect 104990 119200 105046 120000
rect 106554 119200 106610 120000
rect 108118 119200 108174 120000
rect 109682 119200 109738 120000
rect 111246 119200 111302 120000
rect 112810 119200 112866 120000
rect 114466 119200 114522 120000
rect 116030 119200 116086 120000
rect 117594 119200 117650 120000
rect 119158 119200 119214 120000
rect 120722 119200 120778 120000
rect 122286 119200 122342 120000
rect 123942 119200 123998 120000
rect 125506 119200 125562 120000
rect 127070 119200 127126 120000
rect 128634 119200 128690 120000
rect 130198 119200 130254 120000
rect 131762 119200 131818 120000
rect 133418 119200 133474 120000
rect 134982 119200 135038 120000
rect 136546 119200 136602 120000
rect 138110 119200 138166 120000
rect 139674 119200 139730 120000
rect 141238 119200 141294 120000
rect 142894 119200 142950 120000
rect 144458 119200 144514 120000
rect 146022 119200 146078 120000
rect 147586 119200 147642 120000
rect 149150 119200 149206 120000
rect 150714 119200 150770 120000
rect 152370 119200 152426 120000
rect 153934 119200 153990 120000
rect 155498 119200 155554 120000
rect 157062 119200 157118 120000
rect 158626 119200 158682 120000
rect 160190 119200 160246 120000
rect 161846 119200 161902 120000
rect 163410 119200 163466 120000
rect 164974 119200 165030 120000
rect 166538 119200 166594 120000
rect 168102 119200 168158 120000
rect 169666 119200 169722 120000
rect 171322 119200 171378 120000
rect 172886 119200 172942 120000
rect 174450 119200 174506 120000
rect 176014 119200 176070 120000
rect 177578 119200 177634 120000
rect 179142 119200 179198 120000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23202 0 23258 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25410 0 25466 800
rect 25778 0 25834 800
rect 26054 0 26110 800
rect 26422 0 26478 800
rect 26790 0 26846 800
rect 27158 0 27214 800
rect 27526 0 27582 800
rect 27894 0 27950 800
rect 28262 0 28318 800
rect 28630 0 28686 800
rect 28998 0 29054 800
rect 29366 0 29422 800
rect 29734 0 29790 800
rect 30102 0 30158 800
rect 30470 0 30526 800
rect 30838 0 30894 800
rect 31206 0 31262 800
rect 31574 0 31630 800
rect 31942 0 31998 800
rect 32310 0 32366 800
rect 32678 0 32734 800
rect 33046 0 33102 800
rect 33414 0 33470 800
rect 33782 0 33838 800
rect 34150 0 34206 800
rect 34518 0 34574 800
rect 34886 0 34942 800
rect 35254 0 35310 800
rect 35622 0 35678 800
rect 35990 0 36046 800
rect 36358 0 36414 800
rect 36726 0 36782 800
rect 37094 0 37150 800
rect 37462 0 37518 800
rect 37830 0 37886 800
rect 38198 0 38254 800
rect 38566 0 38622 800
rect 38934 0 38990 800
rect 39302 0 39358 800
rect 39670 0 39726 800
rect 40038 0 40094 800
rect 40406 0 40462 800
rect 40774 0 40830 800
rect 41142 0 41198 800
rect 41510 0 41566 800
rect 41878 0 41934 800
rect 42246 0 42302 800
rect 42614 0 42670 800
rect 42982 0 43038 800
rect 43350 0 43406 800
rect 43718 0 43774 800
rect 44086 0 44142 800
rect 44454 0 44510 800
rect 44822 0 44878 800
rect 45190 0 45246 800
rect 45558 0 45614 800
rect 45926 0 45982 800
rect 46294 0 46350 800
rect 46662 0 46718 800
rect 47030 0 47086 800
rect 47398 0 47454 800
rect 47766 0 47822 800
rect 48134 0 48190 800
rect 48502 0 48558 800
rect 48870 0 48926 800
rect 49238 0 49294 800
rect 49606 0 49662 800
rect 49974 0 50030 800
rect 50342 0 50398 800
rect 50710 0 50766 800
rect 51078 0 51134 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 52090 0 52146 800
rect 52458 0 52514 800
rect 52826 0 52882 800
rect 53194 0 53250 800
rect 53562 0 53618 800
rect 53930 0 53986 800
rect 54298 0 54354 800
rect 54666 0 54722 800
rect 55034 0 55090 800
rect 55402 0 55458 800
rect 55770 0 55826 800
rect 56138 0 56194 800
rect 56506 0 56562 800
rect 56874 0 56930 800
rect 57242 0 57298 800
rect 57610 0 57666 800
rect 57978 0 58034 800
rect 58346 0 58402 800
rect 58714 0 58770 800
rect 59082 0 59138 800
rect 59450 0 59506 800
rect 59818 0 59874 800
rect 60186 0 60242 800
rect 60554 0 60610 800
rect 60922 0 60978 800
rect 61290 0 61346 800
rect 61658 0 61714 800
rect 62026 0 62082 800
rect 62394 0 62450 800
rect 62762 0 62818 800
rect 63130 0 63186 800
rect 63498 0 63554 800
rect 63866 0 63922 800
rect 64234 0 64290 800
rect 64602 0 64658 800
rect 64970 0 65026 800
rect 65338 0 65394 800
rect 65706 0 65762 800
rect 66074 0 66130 800
rect 66442 0 66498 800
rect 66810 0 66866 800
rect 67178 0 67234 800
rect 67546 0 67602 800
rect 67914 0 67970 800
rect 68282 0 68338 800
rect 68650 0 68706 800
rect 69018 0 69074 800
rect 69386 0 69442 800
rect 69754 0 69810 800
rect 70122 0 70178 800
rect 70490 0 70546 800
rect 70858 0 70914 800
rect 71226 0 71282 800
rect 71594 0 71650 800
rect 71962 0 72018 800
rect 72330 0 72386 800
rect 72698 0 72754 800
rect 73066 0 73122 800
rect 73434 0 73490 800
rect 73802 0 73858 800
rect 74170 0 74226 800
rect 74538 0 74594 800
rect 74906 0 74962 800
rect 75274 0 75330 800
rect 75642 0 75698 800
rect 76010 0 76066 800
rect 76378 0 76434 800
rect 76746 0 76802 800
rect 77114 0 77170 800
rect 77390 0 77446 800
rect 77758 0 77814 800
rect 78126 0 78182 800
rect 78494 0 78550 800
rect 78862 0 78918 800
rect 79230 0 79286 800
rect 79598 0 79654 800
rect 79966 0 80022 800
rect 80334 0 80390 800
rect 80702 0 80758 800
rect 81070 0 81126 800
rect 81438 0 81494 800
rect 81806 0 81862 800
rect 82174 0 82230 800
rect 82542 0 82598 800
rect 82910 0 82966 800
rect 83278 0 83334 800
rect 83646 0 83702 800
rect 84014 0 84070 800
rect 84382 0 84438 800
rect 84750 0 84806 800
rect 85118 0 85174 800
rect 85486 0 85542 800
rect 85854 0 85910 800
rect 86222 0 86278 800
rect 86590 0 86646 800
rect 86958 0 87014 800
rect 87326 0 87382 800
rect 87694 0 87750 800
rect 88062 0 88118 800
rect 88430 0 88486 800
rect 88798 0 88854 800
rect 89166 0 89222 800
rect 89534 0 89590 800
rect 89902 0 89958 800
rect 90270 0 90326 800
rect 90638 0 90694 800
rect 91006 0 91062 800
rect 91374 0 91430 800
rect 91742 0 91798 800
rect 92110 0 92166 800
rect 92478 0 92534 800
rect 92846 0 92902 800
rect 93214 0 93270 800
rect 93582 0 93638 800
rect 93950 0 94006 800
rect 94318 0 94374 800
rect 94686 0 94742 800
rect 95054 0 95110 800
rect 95422 0 95478 800
rect 95790 0 95846 800
rect 96158 0 96214 800
rect 96526 0 96582 800
rect 96894 0 96950 800
rect 97262 0 97318 800
rect 97630 0 97686 800
rect 97998 0 98054 800
rect 98366 0 98422 800
rect 98734 0 98790 800
rect 99102 0 99158 800
rect 99470 0 99526 800
rect 99838 0 99894 800
rect 100206 0 100262 800
rect 100574 0 100630 800
rect 100942 0 100998 800
rect 101310 0 101366 800
rect 101678 0 101734 800
rect 102046 0 102102 800
rect 102414 0 102470 800
rect 102782 0 102838 800
rect 103058 0 103114 800
rect 103426 0 103482 800
rect 103794 0 103850 800
rect 104162 0 104218 800
rect 104530 0 104586 800
rect 104898 0 104954 800
rect 105266 0 105322 800
rect 105634 0 105690 800
rect 106002 0 106058 800
rect 106370 0 106426 800
rect 106738 0 106794 800
rect 107106 0 107162 800
rect 107474 0 107530 800
rect 107842 0 107898 800
rect 108210 0 108266 800
rect 108578 0 108634 800
rect 108946 0 109002 800
rect 109314 0 109370 800
rect 109682 0 109738 800
rect 110050 0 110106 800
rect 110418 0 110474 800
rect 110786 0 110842 800
rect 111154 0 111210 800
rect 111522 0 111578 800
rect 111890 0 111946 800
rect 112258 0 112314 800
rect 112626 0 112682 800
rect 112994 0 113050 800
rect 113362 0 113418 800
rect 113730 0 113786 800
rect 114098 0 114154 800
rect 114466 0 114522 800
rect 114834 0 114890 800
rect 115202 0 115258 800
rect 115570 0 115626 800
rect 115938 0 115994 800
rect 116306 0 116362 800
rect 116674 0 116730 800
rect 117042 0 117098 800
rect 117410 0 117466 800
rect 117778 0 117834 800
rect 118146 0 118202 800
rect 118514 0 118570 800
rect 118882 0 118938 800
rect 119250 0 119306 800
rect 119618 0 119674 800
rect 119986 0 120042 800
rect 120354 0 120410 800
rect 120722 0 120778 800
rect 121090 0 121146 800
rect 121458 0 121514 800
rect 121826 0 121882 800
rect 122194 0 122250 800
rect 122562 0 122618 800
rect 122930 0 122986 800
rect 123298 0 123354 800
rect 123666 0 123722 800
rect 124034 0 124090 800
rect 124402 0 124458 800
rect 124770 0 124826 800
rect 125138 0 125194 800
rect 125506 0 125562 800
rect 125874 0 125930 800
rect 126242 0 126298 800
rect 126610 0 126666 800
rect 126978 0 127034 800
rect 127346 0 127402 800
rect 127714 0 127770 800
rect 128082 0 128138 800
rect 128450 0 128506 800
rect 128726 0 128782 800
rect 129094 0 129150 800
rect 129462 0 129518 800
rect 129830 0 129886 800
rect 130198 0 130254 800
rect 130566 0 130622 800
rect 130934 0 130990 800
rect 131302 0 131358 800
rect 131670 0 131726 800
rect 132038 0 132094 800
rect 132406 0 132462 800
rect 132774 0 132830 800
rect 133142 0 133198 800
rect 133510 0 133566 800
rect 133878 0 133934 800
rect 134246 0 134302 800
rect 134614 0 134670 800
rect 134982 0 135038 800
rect 135350 0 135406 800
rect 135718 0 135774 800
rect 136086 0 136142 800
rect 136454 0 136510 800
rect 136822 0 136878 800
rect 137190 0 137246 800
rect 137558 0 137614 800
rect 137926 0 137982 800
rect 138294 0 138350 800
rect 138662 0 138718 800
rect 139030 0 139086 800
rect 139398 0 139454 800
rect 139766 0 139822 800
rect 140134 0 140190 800
rect 140502 0 140558 800
rect 140870 0 140926 800
rect 141238 0 141294 800
rect 141606 0 141662 800
rect 141974 0 142030 800
rect 142342 0 142398 800
rect 142710 0 142766 800
rect 143078 0 143134 800
rect 143446 0 143502 800
rect 143814 0 143870 800
rect 144182 0 144238 800
rect 144550 0 144606 800
rect 144918 0 144974 800
rect 145286 0 145342 800
rect 145654 0 145710 800
rect 146022 0 146078 800
rect 146390 0 146446 800
rect 146758 0 146814 800
rect 147126 0 147182 800
rect 147494 0 147550 800
rect 147862 0 147918 800
rect 148230 0 148286 800
rect 148598 0 148654 800
rect 148966 0 149022 800
rect 149334 0 149390 800
rect 149702 0 149758 800
rect 150070 0 150126 800
rect 150438 0 150494 800
rect 150806 0 150862 800
rect 151174 0 151230 800
rect 151542 0 151598 800
rect 151910 0 151966 800
rect 152278 0 152334 800
rect 152646 0 152702 800
rect 153014 0 153070 800
rect 153382 0 153438 800
rect 153750 0 153806 800
rect 154118 0 154174 800
rect 154394 0 154450 800
rect 154762 0 154818 800
rect 155130 0 155186 800
rect 155498 0 155554 800
rect 155866 0 155922 800
rect 156234 0 156290 800
rect 156602 0 156658 800
rect 156970 0 157026 800
rect 157338 0 157394 800
rect 157706 0 157762 800
rect 158074 0 158130 800
rect 158442 0 158498 800
rect 158810 0 158866 800
rect 159178 0 159234 800
rect 159546 0 159602 800
rect 159914 0 159970 800
rect 160282 0 160338 800
rect 160650 0 160706 800
rect 161018 0 161074 800
rect 161386 0 161442 800
rect 161754 0 161810 800
rect 162122 0 162178 800
rect 162490 0 162546 800
rect 162858 0 162914 800
rect 163226 0 163282 800
rect 163594 0 163650 800
rect 163962 0 164018 800
rect 164330 0 164386 800
rect 164698 0 164754 800
rect 165066 0 165122 800
rect 165434 0 165490 800
rect 165802 0 165858 800
rect 166170 0 166226 800
rect 166538 0 166594 800
rect 166906 0 166962 800
rect 167274 0 167330 800
rect 167642 0 167698 800
rect 168010 0 168066 800
rect 168378 0 168434 800
rect 168746 0 168802 800
rect 169114 0 169170 800
rect 169482 0 169538 800
rect 169850 0 169906 800
rect 170218 0 170274 800
rect 170586 0 170642 800
rect 170954 0 171010 800
rect 171322 0 171378 800
rect 171690 0 171746 800
rect 172058 0 172114 800
rect 172426 0 172482 800
rect 172794 0 172850 800
rect 173162 0 173218 800
rect 173530 0 173586 800
rect 173898 0 173954 800
rect 174266 0 174322 800
rect 174634 0 174690 800
rect 175002 0 175058 800
rect 175370 0 175426 800
rect 175738 0 175794 800
rect 176106 0 176162 800
rect 176474 0 176530 800
rect 176842 0 176898 800
rect 177210 0 177266 800
rect 177578 0 177634 800
rect 177946 0 178002 800
rect 178314 0 178370 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
<< obsm2 >>
rect 112 119144 698 119200
rect 866 119144 2262 119200
rect 2430 119144 3826 119200
rect 3994 119144 5390 119200
rect 5558 119144 6954 119200
rect 7122 119144 8518 119200
rect 8686 119144 10174 119200
rect 10342 119144 11738 119200
rect 11906 119144 13302 119200
rect 13470 119144 14866 119200
rect 15034 119144 16430 119200
rect 16598 119144 17994 119200
rect 18162 119144 19650 119200
rect 19818 119144 21214 119200
rect 21382 119144 22778 119200
rect 22946 119144 24342 119200
rect 24510 119144 25906 119200
rect 26074 119144 27470 119200
rect 27638 119144 29126 119200
rect 29294 119144 30690 119200
rect 30858 119144 32254 119200
rect 32422 119144 33818 119200
rect 33986 119144 35382 119200
rect 35550 119144 36946 119200
rect 37114 119144 38602 119200
rect 38770 119144 40166 119200
rect 40334 119144 41730 119200
rect 41898 119144 43294 119200
rect 43462 119144 44858 119200
rect 45026 119144 46422 119200
rect 46590 119144 48078 119200
rect 48246 119144 49642 119200
rect 49810 119144 51206 119200
rect 51374 119144 52770 119200
rect 52938 119144 54334 119200
rect 54502 119144 55898 119200
rect 56066 119144 57554 119200
rect 57722 119144 59118 119200
rect 59286 119144 60682 119200
rect 60850 119144 62246 119200
rect 62414 119144 63810 119200
rect 63978 119144 65374 119200
rect 65542 119144 67030 119200
rect 67198 119144 68594 119200
rect 68762 119144 70158 119200
rect 70326 119144 71722 119200
rect 71890 119144 73286 119200
rect 73454 119144 74850 119200
rect 75018 119144 76506 119200
rect 76674 119144 78070 119200
rect 78238 119144 79634 119200
rect 79802 119144 81198 119200
rect 81366 119144 82762 119200
rect 82930 119144 84326 119200
rect 84494 119144 85982 119200
rect 86150 119144 87546 119200
rect 87714 119144 89110 119200
rect 89278 119144 90674 119200
rect 90842 119144 92238 119200
rect 92406 119144 93802 119200
rect 93970 119144 95458 119200
rect 95626 119144 97022 119200
rect 97190 119144 98586 119200
rect 98754 119144 100150 119200
rect 100318 119144 101714 119200
rect 101882 119144 103278 119200
rect 103446 119144 104934 119200
rect 105102 119144 106498 119200
rect 106666 119144 108062 119200
rect 108230 119144 109626 119200
rect 109794 119144 111190 119200
rect 111358 119144 112754 119200
rect 112922 119144 114410 119200
rect 114578 119144 115974 119200
rect 116142 119144 117538 119200
rect 117706 119144 119102 119200
rect 119270 119144 120666 119200
rect 120834 119144 122230 119200
rect 122398 119144 123886 119200
rect 124054 119144 125450 119200
rect 125618 119144 127014 119200
rect 127182 119144 128578 119200
rect 128746 119144 130142 119200
rect 130310 119144 131706 119200
rect 131874 119144 133362 119200
rect 133530 119144 134926 119200
rect 135094 119144 136490 119200
rect 136658 119144 138054 119200
rect 138222 119144 139618 119200
rect 139786 119144 141182 119200
rect 141350 119144 142838 119200
rect 143006 119144 144402 119200
rect 144570 119144 145966 119200
rect 146134 119144 147530 119200
rect 147698 119144 149094 119200
rect 149262 119144 150658 119200
rect 150826 119144 152314 119200
rect 152482 119144 153878 119200
rect 154046 119144 155442 119200
rect 155610 119144 157006 119200
rect 157174 119144 158570 119200
rect 158738 119144 160134 119200
rect 160302 119144 161790 119200
rect 161958 119144 163354 119200
rect 163522 119144 164918 119200
rect 165086 119144 166482 119200
rect 166650 119144 168046 119200
rect 168214 119144 169610 119200
rect 169778 119144 171266 119200
rect 171434 119144 172830 119200
rect 172998 119144 174394 119200
rect 174562 119144 175958 119200
rect 176126 119144 177522 119200
rect 177690 119144 179086 119200
rect 179254 119144 179840 119200
rect 112 856 179840 119144
rect 222 342 330 856
rect 498 342 698 856
rect 866 342 1066 856
rect 1234 342 1434 856
rect 1602 342 1802 856
rect 1970 342 2170 856
rect 2338 342 2538 856
rect 2706 342 2906 856
rect 3074 342 3274 856
rect 3442 342 3642 856
rect 3810 342 4010 856
rect 4178 342 4378 856
rect 4546 342 4746 856
rect 4914 342 5114 856
rect 5282 342 5482 856
rect 5650 342 5850 856
rect 6018 342 6218 856
rect 6386 342 6586 856
rect 6754 342 6954 856
rect 7122 342 7322 856
rect 7490 342 7690 856
rect 7858 342 8058 856
rect 8226 342 8426 856
rect 8594 342 8794 856
rect 8962 342 9162 856
rect 9330 342 9530 856
rect 9698 342 9898 856
rect 10066 342 10266 856
rect 10434 342 10634 856
rect 10802 342 11002 856
rect 11170 342 11370 856
rect 11538 342 11738 856
rect 11906 342 12106 856
rect 12274 342 12474 856
rect 12642 342 12842 856
rect 13010 342 13210 856
rect 13378 342 13578 856
rect 13746 342 13946 856
rect 14114 342 14314 856
rect 14482 342 14682 856
rect 14850 342 15050 856
rect 15218 342 15418 856
rect 15586 342 15786 856
rect 15954 342 16154 856
rect 16322 342 16522 856
rect 16690 342 16890 856
rect 17058 342 17258 856
rect 17426 342 17626 856
rect 17794 342 17994 856
rect 18162 342 18362 856
rect 18530 342 18730 856
rect 18898 342 19098 856
rect 19266 342 19466 856
rect 19634 342 19834 856
rect 20002 342 20202 856
rect 20370 342 20570 856
rect 20738 342 20938 856
rect 21106 342 21306 856
rect 21474 342 21674 856
rect 21842 342 22042 856
rect 22210 342 22410 856
rect 22578 342 22778 856
rect 22946 342 23146 856
rect 23314 342 23514 856
rect 23682 342 23882 856
rect 24050 342 24250 856
rect 24418 342 24618 856
rect 24786 342 24986 856
rect 25154 342 25354 856
rect 25522 342 25722 856
rect 25890 342 25998 856
rect 26166 342 26366 856
rect 26534 342 26734 856
rect 26902 342 27102 856
rect 27270 342 27470 856
rect 27638 342 27838 856
rect 28006 342 28206 856
rect 28374 342 28574 856
rect 28742 342 28942 856
rect 29110 342 29310 856
rect 29478 342 29678 856
rect 29846 342 30046 856
rect 30214 342 30414 856
rect 30582 342 30782 856
rect 30950 342 31150 856
rect 31318 342 31518 856
rect 31686 342 31886 856
rect 32054 342 32254 856
rect 32422 342 32622 856
rect 32790 342 32990 856
rect 33158 342 33358 856
rect 33526 342 33726 856
rect 33894 342 34094 856
rect 34262 342 34462 856
rect 34630 342 34830 856
rect 34998 342 35198 856
rect 35366 342 35566 856
rect 35734 342 35934 856
rect 36102 342 36302 856
rect 36470 342 36670 856
rect 36838 342 37038 856
rect 37206 342 37406 856
rect 37574 342 37774 856
rect 37942 342 38142 856
rect 38310 342 38510 856
rect 38678 342 38878 856
rect 39046 342 39246 856
rect 39414 342 39614 856
rect 39782 342 39982 856
rect 40150 342 40350 856
rect 40518 342 40718 856
rect 40886 342 41086 856
rect 41254 342 41454 856
rect 41622 342 41822 856
rect 41990 342 42190 856
rect 42358 342 42558 856
rect 42726 342 42926 856
rect 43094 342 43294 856
rect 43462 342 43662 856
rect 43830 342 44030 856
rect 44198 342 44398 856
rect 44566 342 44766 856
rect 44934 342 45134 856
rect 45302 342 45502 856
rect 45670 342 45870 856
rect 46038 342 46238 856
rect 46406 342 46606 856
rect 46774 342 46974 856
rect 47142 342 47342 856
rect 47510 342 47710 856
rect 47878 342 48078 856
rect 48246 342 48446 856
rect 48614 342 48814 856
rect 48982 342 49182 856
rect 49350 342 49550 856
rect 49718 342 49918 856
rect 50086 342 50286 856
rect 50454 342 50654 856
rect 50822 342 51022 856
rect 51190 342 51390 856
rect 51558 342 51666 856
rect 51834 342 52034 856
rect 52202 342 52402 856
rect 52570 342 52770 856
rect 52938 342 53138 856
rect 53306 342 53506 856
rect 53674 342 53874 856
rect 54042 342 54242 856
rect 54410 342 54610 856
rect 54778 342 54978 856
rect 55146 342 55346 856
rect 55514 342 55714 856
rect 55882 342 56082 856
rect 56250 342 56450 856
rect 56618 342 56818 856
rect 56986 342 57186 856
rect 57354 342 57554 856
rect 57722 342 57922 856
rect 58090 342 58290 856
rect 58458 342 58658 856
rect 58826 342 59026 856
rect 59194 342 59394 856
rect 59562 342 59762 856
rect 59930 342 60130 856
rect 60298 342 60498 856
rect 60666 342 60866 856
rect 61034 342 61234 856
rect 61402 342 61602 856
rect 61770 342 61970 856
rect 62138 342 62338 856
rect 62506 342 62706 856
rect 62874 342 63074 856
rect 63242 342 63442 856
rect 63610 342 63810 856
rect 63978 342 64178 856
rect 64346 342 64546 856
rect 64714 342 64914 856
rect 65082 342 65282 856
rect 65450 342 65650 856
rect 65818 342 66018 856
rect 66186 342 66386 856
rect 66554 342 66754 856
rect 66922 342 67122 856
rect 67290 342 67490 856
rect 67658 342 67858 856
rect 68026 342 68226 856
rect 68394 342 68594 856
rect 68762 342 68962 856
rect 69130 342 69330 856
rect 69498 342 69698 856
rect 69866 342 70066 856
rect 70234 342 70434 856
rect 70602 342 70802 856
rect 70970 342 71170 856
rect 71338 342 71538 856
rect 71706 342 71906 856
rect 72074 342 72274 856
rect 72442 342 72642 856
rect 72810 342 73010 856
rect 73178 342 73378 856
rect 73546 342 73746 856
rect 73914 342 74114 856
rect 74282 342 74482 856
rect 74650 342 74850 856
rect 75018 342 75218 856
rect 75386 342 75586 856
rect 75754 342 75954 856
rect 76122 342 76322 856
rect 76490 342 76690 856
rect 76858 342 77058 856
rect 77226 342 77334 856
rect 77502 342 77702 856
rect 77870 342 78070 856
rect 78238 342 78438 856
rect 78606 342 78806 856
rect 78974 342 79174 856
rect 79342 342 79542 856
rect 79710 342 79910 856
rect 80078 342 80278 856
rect 80446 342 80646 856
rect 80814 342 81014 856
rect 81182 342 81382 856
rect 81550 342 81750 856
rect 81918 342 82118 856
rect 82286 342 82486 856
rect 82654 342 82854 856
rect 83022 342 83222 856
rect 83390 342 83590 856
rect 83758 342 83958 856
rect 84126 342 84326 856
rect 84494 342 84694 856
rect 84862 342 85062 856
rect 85230 342 85430 856
rect 85598 342 85798 856
rect 85966 342 86166 856
rect 86334 342 86534 856
rect 86702 342 86902 856
rect 87070 342 87270 856
rect 87438 342 87638 856
rect 87806 342 88006 856
rect 88174 342 88374 856
rect 88542 342 88742 856
rect 88910 342 89110 856
rect 89278 342 89478 856
rect 89646 342 89846 856
rect 90014 342 90214 856
rect 90382 342 90582 856
rect 90750 342 90950 856
rect 91118 342 91318 856
rect 91486 342 91686 856
rect 91854 342 92054 856
rect 92222 342 92422 856
rect 92590 342 92790 856
rect 92958 342 93158 856
rect 93326 342 93526 856
rect 93694 342 93894 856
rect 94062 342 94262 856
rect 94430 342 94630 856
rect 94798 342 94998 856
rect 95166 342 95366 856
rect 95534 342 95734 856
rect 95902 342 96102 856
rect 96270 342 96470 856
rect 96638 342 96838 856
rect 97006 342 97206 856
rect 97374 342 97574 856
rect 97742 342 97942 856
rect 98110 342 98310 856
rect 98478 342 98678 856
rect 98846 342 99046 856
rect 99214 342 99414 856
rect 99582 342 99782 856
rect 99950 342 100150 856
rect 100318 342 100518 856
rect 100686 342 100886 856
rect 101054 342 101254 856
rect 101422 342 101622 856
rect 101790 342 101990 856
rect 102158 342 102358 856
rect 102526 342 102726 856
rect 102894 342 103002 856
rect 103170 342 103370 856
rect 103538 342 103738 856
rect 103906 342 104106 856
rect 104274 342 104474 856
rect 104642 342 104842 856
rect 105010 342 105210 856
rect 105378 342 105578 856
rect 105746 342 105946 856
rect 106114 342 106314 856
rect 106482 342 106682 856
rect 106850 342 107050 856
rect 107218 342 107418 856
rect 107586 342 107786 856
rect 107954 342 108154 856
rect 108322 342 108522 856
rect 108690 342 108890 856
rect 109058 342 109258 856
rect 109426 342 109626 856
rect 109794 342 109994 856
rect 110162 342 110362 856
rect 110530 342 110730 856
rect 110898 342 111098 856
rect 111266 342 111466 856
rect 111634 342 111834 856
rect 112002 342 112202 856
rect 112370 342 112570 856
rect 112738 342 112938 856
rect 113106 342 113306 856
rect 113474 342 113674 856
rect 113842 342 114042 856
rect 114210 342 114410 856
rect 114578 342 114778 856
rect 114946 342 115146 856
rect 115314 342 115514 856
rect 115682 342 115882 856
rect 116050 342 116250 856
rect 116418 342 116618 856
rect 116786 342 116986 856
rect 117154 342 117354 856
rect 117522 342 117722 856
rect 117890 342 118090 856
rect 118258 342 118458 856
rect 118626 342 118826 856
rect 118994 342 119194 856
rect 119362 342 119562 856
rect 119730 342 119930 856
rect 120098 342 120298 856
rect 120466 342 120666 856
rect 120834 342 121034 856
rect 121202 342 121402 856
rect 121570 342 121770 856
rect 121938 342 122138 856
rect 122306 342 122506 856
rect 122674 342 122874 856
rect 123042 342 123242 856
rect 123410 342 123610 856
rect 123778 342 123978 856
rect 124146 342 124346 856
rect 124514 342 124714 856
rect 124882 342 125082 856
rect 125250 342 125450 856
rect 125618 342 125818 856
rect 125986 342 126186 856
rect 126354 342 126554 856
rect 126722 342 126922 856
rect 127090 342 127290 856
rect 127458 342 127658 856
rect 127826 342 128026 856
rect 128194 342 128394 856
rect 128562 342 128670 856
rect 128838 342 129038 856
rect 129206 342 129406 856
rect 129574 342 129774 856
rect 129942 342 130142 856
rect 130310 342 130510 856
rect 130678 342 130878 856
rect 131046 342 131246 856
rect 131414 342 131614 856
rect 131782 342 131982 856
rect 132150 342 132350 856
rect 132518 342 132718 856
rect 132886 342 133086 856
rect 133254 342 133454 856
rect 133622 342 133822 856
rect 133990 342 134190 856
rect 134358 342 134558 856
rect 134726 342 134926 856
rect 135094 342 135294 856
rect 135462 342 135662 856
rect 135830 342 136030 856
rect 136198 342 136398 856
rect 136566 342 136766 856
rect 136934 342 137134 856
rect 137302 342 137502 856
rect 137670 342 137870 856
rect 138038 342 138238 856
rect 138406 342 138606 856
rect 138774 342 138974 856
rect 139142 342 139342 856
rect 139510 342 139710 856
rect 139878 342 140078 856
rect 140246 342 140446 856
rect 140614 342 140814 856
rect 140982 342 141182 856
rect 141350 342 141550 856
rect 141718 342 141918 856
rect 142086 342 142286 856
rect 142454 342 142654 856
rect 142822 342 143022 856
rect 143190 342 143390 856
rect 143558 342 143758 856
rect 143926 342 144126 856
rect 144294 342 144494 856
rect 144662 342 144862 856
rect 145030 342 145230 856
rect 145398 342 145598 856
rect 145766 342 145966 856
rect 146134 342 146334 856
rect 146502 342 146702 856
rect 146870 342 147070 856
rect 147238 342 147438 856
rect 147606 342 147806 856
rect 147974 342 148174 856
rect 148342 342 148542 856
rect 148710 342 148910 856
rect 149078 342 149278 856
rect 149446 342 149646 856
rect 149814 342 150014 856
rect 150182 342 150382 856
rect 150550 342 150750 856
rect 150918 342 151118 856
rect 151286 342 151486 856
rect 151654 342 151854 856
rect 152022 342 152222 856
rect 152390 342 152590 856
rect 152758 342 152958 856
rect 153126 342 153326 856
rect 153494 342 153694 856
rect 153862 342 154062 856
rect 154230 342 154338 856
rect 154506 342 154706 856
rect 154874 342 155074 856
rect 155242 342 155442 856
rect 155610 342 155810 856
rect 155978 342 156178 856
rect 156346 342 156546 856
rect 156714 342 156914 856
rect 157082 342 157282 856
rect 157450 342 157650 856
rect 157818 342 158018 856
rect 158186 342 158386 856
rect 158554 342 158754 856
rect 158922 342 159122 856
rect 159290 342 159490 856
rect 159658 342 159858 856
rect 160026 342 160226 856
rect 160394 342 160594 856
rect 160762 342 160962 856
rect 161130 342 161330 856
rect 161498 342 161698 856
rect 161866 342 162066 856
rect 162234 342 162434 856
rect 162602 342 162802 856
rect 162970 342 163170 856
rect 163338 342 163538 856
rect 163706 342 163906 856
rect 164074 342 164274 856
rect 164442 342 164642 856
rect 164810 342 165010 856
rect 165178 342 165378 856
rect 165546 342 165746 856
rect 165914 342 166114 856
rect 166282 342 166482 856
rect 166650 342 166850 856
rect 167018 342 167218 856
rect 167386 342 167586 856
rect 167754 342 167954 856
rect 168122 342 168322 856
rect 168490 342 168690 856
rect 168858 342 169058 856
rect 169226 342 169426 856
rect 169594 342 169794 856
rect 169962 342 170162 856
rect 170330 342 170530 856
rect 170698 342 170898 856
rect 171066 342 171266 856
rect 171434 342 171634 856
rect 171802 342 172002 856
rect 172170 342 172370 856
rect 172538 342 172738 856
rect 172906 342 173106 856
rect 173274 342 173474 856
rect 173642 342 173842 856
rect 174010 342 174210 856
rect 174378 342 174578 856
rect 174746 342 174946 856
rect 175114 342 175314 856
rect 175482 342 175682 856
rect 175850 342 176050 856
rect 176218 342 176418 856
rect 176586 342 176786 856
rect 176954 342 177154 856
rect 177322 342 177522 856
rect 177690 342 177890 856
rect 178058 342 178258 856
rect 178426 342 178626 856
rect 178794 342 178994 856
rect 179162 342 179362 856
rect 179530 342 179730 856
<< metal3 >>
rect 0 89904 800 90024
rect 0 29928 800 30048
<< obsm3 >>
rect 800 90104 173488 117537
rect 880 89824 173488 90104
rect 800 30128 173488 89824
rect 880 29848 173488 30128
rect 800 1803 173488 29848
<< metal4 >>
rect 4208 2128 4528 117552
rect 4868 2176 5188 117504
rect 5528 2176 5848 117504
rect 6188 2176 6508 117504
rect 19568 2128 19888 117552
rect 20228 2176 20548 117504
rect 20888 2176 21208 117504
rect 21548 2176 21868 117504
rect 34928 2128 35248 117552
rect 35588 2176 35908 117504
rect 36248 2176 36568 117504
rect 36908 2176 37228 117504
rect 50288 2128 50608 117552
rect 50948 2176 51268 117504
rect 51608 2176 51928 117504
rect 52268 2176 52588 117504
rect 65648 2128 65968 117552
rect 66308 2176 66628 117504
rect 66968 2176 67288 117504
rect 67628 2176 67948 117504
rect 81008 2128 81328 117552
rect 81668 2176 81988 117504
rect 82328 2176 82648 117504
rect 82988 2176 83308 117504
rect 96368 2128 96688 117552
rect 97028 2176 97348 117504
rect 97688 2176 98008 117504
rect 98348 2176 98668 117504
rect 111728 2128 112048 117552
rect 112388 2176 112708 117504
rect 113048 2176 113368 117504
rect 113708 2176 114028 117504
rect 127088 2128 127408 117552
rect 127748 2176 128068 117504
rect 128408 2176 128728 117504
rect 129068 2176 129388 117504
rect 142448 2128 142768 117552
rect 143108 2176 143428 117504
rect 143768 2176 144088 117504
rect 144428 2176 144748 117504
rect 157808 2128 158128 117552
rect 158468 2176 158788 117504
rect 159128 2176 159448 117504
rect 159788 2176 160108 117504
rect 173168 2128 173488 117552
rect 173828 2176 174148 117504
rect 174488 2176 174808 117504
rect 175148 2176 175468 117504
<< obsm4 >>
rect 2550 2075 4128 6629
rect 4608 2096 4788 6629
rect 5268 2096 5448 6629
rect 5928 2096 6108 6629
rect 6588 2096 19488 6629
rect 4608 2075 19488 2096
rect 19968 2096 20148 6629
rect 20628 2096 20808 6629
rect 21288 2096 21468 6629
rect 21948 2096 34848 6629
rect 19968 2075 34848 2096
rect 35328 2096 35508 6629
rect 35988 2096 36168 6629
rect 36648 2096 36828 6629
rect 37308 2096 50208 6629
rect 35328 2075 50208 2096
rect 50688 2096 50868 6629
rect 51348 2096 51528 6629
rect 52008 2096 52188 6629
rect 52668 2096 65568 6629
rect 50688 2075 65568 2096
rect 66048 2096 66228 6629
rect 66708 2096 66888 6629
rect 67368 2096 67548 6629
rect 68028 2096 80928 6629
rect 66048 2075 80928 2096
rect 81408 2096 81588 6629
rect 82068 2096 82248 6629
rect 82728 2096 82908 6629
rect 83388 2096 96288 6629
rect 81408 2075 96288 2096
rect 96768 2096 96948 6629
rect 97428 2096 97608 6629
rect 98088 2096 98268 6629
rect 98748 2096 100858 6629
rect 96768 2075 100858 2096
<< obsm5 >>
rect 2508 2900 100900 3220
<< labels >>
rlabel metal2 s 754 119200 810 120000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 48134 119200 48190 120000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 52826 119200 52882 120000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 57610 119200 57666 120000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 62302 119200 62358 120000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 67086 119200 67142 120000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 71778 119200 71834 120000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 76562 119200 76618 120000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 81254 119200 81310 120000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 86038 119200 86094 120000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 90730 119200 90786 120000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 5446 119200 5502 120000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 95514 119200 95570 120000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 100206 119200 100262 120000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 104990 119200 105046 120000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 109682 119200 109738 120000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 114466 119200 114522 120000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 119158 119200 119214 120000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 123942 119200 123998 120000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 128634 119200 128690 120000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 133418 119200 133474 120000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 138110 119200 138166 120000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 10230 119200 10286 120000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 142894 119200 142950 120000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 147586 119200 147642 120000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 152370 119200 152426 120000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 157062 119200 157118 120000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 161846 119200 161902 120000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 166538 119200 166594 120000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 171322 119200 171378 120000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 176014 119200 176070 120000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 14922 119200 14978 120000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 19706 119200 19762 120000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 24398 119200 24454 120000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 29182 119200 29238 120000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 33874 119200 33930 120000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 38658 119200 38714 120000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 43350 119200 43406 120000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2318 119200 2374 120000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 49698 119200 49754 120000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 54390 119200 54446 120000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 59174 119200 59230 120000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 63866 119200 63922 120000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 68650 119200 68706 120000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 73342 119200 73398 120000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 78126 119200 78182 120000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 82818 119200 82874 120000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 87602 119200 87658 120000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 92294 119200 92350 120000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7010 119200 7066 120000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 97078 119200 97134 120000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 101770 119200 101826 120000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 106554 119200 106610 120000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 111246 119200 111302 120000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 116030 119200 116086 120000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 120722 119200 120778 120000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 125506 119200 125562 120000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 130198 119200 130254 120000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 134982 119200 135038 120000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 139674 119200 139730 120000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 11794 119200 11850 120000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 144458 119200 144514 120000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 149150 119200 149206 120000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 153934 119200 153990 120000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 158626 119200 158682 120000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 163410 119200 163466 120000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 168102 119200 168158 120000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 172886 119200 172942 120000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 177578 119200 177634 120000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 16486 119200 16542 120000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 21270 119200 21326 120000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 25962 119200 26018 120000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 30746 119200 30802 120000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 35438 119200 35494 120000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 40222 119200 40278 120000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 44914 119200 44970 120000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 3882 119200 3938 120000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 51262 119200 51318 120000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 55954 119200 56010 120000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 60738 119200 60794 120000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 65430 119200 65486 120000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 70214 119200 70270 120000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 74906 119200 74962 120000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 79690 119200 79746 120000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 84382 119200 84438 120000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 89166 119200 89222 120000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 93858 119200 93914 120000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 8574 119200 8630 120000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 98642 119200 98698 120000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 103334 119200 103390 120000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 108118 119200 108174 120000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 112810 119200 112866 120000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 117594 119200 117650 120000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 122286 119200 122342 120000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 127070 119200 127126 120000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 131762 119200 131818 120000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 136546 119200 136602 120000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 141238 119200 141294 120000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 13358 119200 13414 120000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 146022 119200 146078 120000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 150714 119200 150770 120000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 155498 119200 155554 120000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 160190 119200 160246 120000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 164974 119200 165030 120000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 169666 119200 169722 120000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 174450 119200 174506 120000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 179142 119200 179198 120000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 18050 119200 18106 120000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 22834 119200 22890 120000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 27526 119200 27582 120000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 32310 119200 32366 120000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 37002 119200 37058 120000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 41786 119200 41842 120000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 46478 119200 46534 120000 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 0 89904 800 90024 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 179786 0 179842 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 148966 0 149022 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 150070 0 150126 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 152278 0 152334 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 153382 0 153438 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 154394 0 154450 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 157706 0 157762 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 158810 0 158866 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 163226 0 163282 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 164330 0 164386 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 165434 0 165490 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 166538 0 166594 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 167642 0 167698 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 168746 0 168802 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 169850 0 169906 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 175370 0 175426 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 177578 0 177634 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 109314 0 109370 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 112626 0 112682 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 120354 0 120410 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 122562 0 122618 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 125874 0 125930 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 129094 0 129150 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 132406 0 132462 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 135718 0 135774 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 139030 0 139086 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 140134 0 140190 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 143446 0 143502 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 144550 0 144606 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 145654 0 145710 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 146758 0 146814 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 147862 0 147918 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 149334 0 149390 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 150438 0 150494 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 151542 0 151598 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 152646 0 152702 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 153750 0 153806 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 154762 0 154818 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 156970 0 157026 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 158074 0 158130 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 159178 0 159234 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 160282 0 160338 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 161386 0 161442 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 162490 0 162546 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 163594 0 163650 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 164698 0 164754 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 165802 0 165858 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 166906 0 166962 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 168010 0 168066 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 169114 0 169170 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 170218 0 170274 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 51446 0 51502 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 171322 0 171378 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 172426 0 172482 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 173530 0 173586 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 174634 0 174690 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 175738 0 175794 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 176842 0 176898 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 177946 0 178002 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 179050 0 179106 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 53562 0 53618 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 61290 0 61346 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 63498 0 63554 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 64602 0 64658 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 70122 0 70178 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 71226 0 71282 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 72330 0 72386 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 76746 0 76802 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 78862 0 78918 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 79966 0 80022 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 82174 0 82230 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 83278 0 83334 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 85486 0 85542 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 86590 0 86646 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 88798 0 88854 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 93214 0 93270 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 95422 0 95478 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 96526 0 96582 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 97630 0 97686 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 98734 0 98790 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 100942 0 100998 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 102046 0 102102 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 103058 0 103114 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 104162 0 104218 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 105266 0 105322 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 106370 0 106426 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 107474 0 107530 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 108578 0 108634 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 109682 0 109738 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 111890 0 111946 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 114098 0 114154 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 115202 0 115258 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 116306 0 116362 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 117410 0 117466 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 119618 0 119674 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 120722 0 120778 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 121826 0 121882 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 122930 0 122986 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 124034 0 124090 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 125138 0 125194 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 126242 0 126298 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 127346 0 127402 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 128450 0 128506 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 129462 0 129518 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 130566 0 130622 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 131670 0 131726 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 132774 0 132830 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 133878 0 133934 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 134982 0 135038 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 136086 0 136142 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 137190 0 137246 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 138294 0 138350 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 139398 0 139454 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 140502 0 140558 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 141606 0 141662 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 142710 0 142766 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 143814 0 143870 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 146022 0 146078 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 147126 0 147182 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 148230 0 148286 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 149702 0 149758 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 150806 0 150862 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 153014 0 153070 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 154118 0 154174 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 155130 0 155186 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 157338 0 157394 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 158442 0 158498 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 159546 0 159602 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 160650 0 160706 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 161754 0 161810 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 162858 0 162914 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 163962 0 164018 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 167274 0 167330 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 168378 0 168434 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 169482 0 169538 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 170586 0 170642 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 171690 0 171746 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 172794 0 172850 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 173898 0 173954 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 175002 0 175058 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 177210 0 177266 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 178314 0 178370 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 179418 0 179474 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 111154 0 111210 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 112258 0 112314 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 114466 0 114522 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 116674 0 116730 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 119986 0 120042 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 122194 0 122250 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 123298 0 123354 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 129830 0 129886 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 130934 0 130990 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 138662 0 138718 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 139766 0 139822 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 141974 0 142030 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 145286 0 145342 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 148598 0 148654 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 504 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[0]
port 570 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_o[10]
port 571 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 wbs_dat_o[11]
port 572 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_o[12]
port 573 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_o[13]
port 574 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 wbs_dat_o[14]
port 575 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_o[15]
port 576 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_o[16]
port 577 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_o[17]
port 578 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_o[18]
port 579 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_o[19]
port 580 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[1]
port 581 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_o[20]
port 582 nsew signal output
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_o[21]
port 583 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_o[22]
port 584 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 wbs_dat_o[23]
port 585 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 wbs_dat_o[24]
port 586 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 wbs_dat_o[25]
port 587 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 wbs_dat_o[26]
port 588 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 wbs_dat_o[27]
port 589 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_o[28]
port 590 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 wbs_dat_o[29]
port 591 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[2]
port 592 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_o[30]
port 593 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 wbs_dat_o[31]
port 594 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[3]
port 595 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_o[4]
port 596 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[5]
port 597 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[6]
port 598 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 wbs_dat_o[7]
port 599 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_o[8]
port 600 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_o[9]
port 601 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_we_i
port 607 nsew signal input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 613 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 614 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 615 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 616 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 617 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 618 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 619 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 117504 6 vccd2
port 620 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 117504 6 vccd2
port 621 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 117504 6 vccd2
port 622 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 117504 6 vccd2
port 623 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 117504 6 vccd2
port 624 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 117504 6 vccd2
port 625 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 117504 6 vssd2
port 626 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 117504 6 vssd2
port 627 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 117504 6 vssd2
port 628 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 117504 6 vssd2
port 629 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 117504 6 vssd2
port 630 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 117504 6 vssd2
port 631 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 117504 6 vdda1
port 632 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 117504 6 vdda1
port 633 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 117504 6 vdda1
port 634 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 117504 6 vdda1
port 635 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 117504 6 vdda1
port 636 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 117504 6 vdda1
port 637 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 117504 6 vssa1
port 638 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 117504 6 vssa1
port 639 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 117504 6 vssa1
port 640 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 117504 6 vssa1
port 641 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 117504 6 vssa1
port 642 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 117504 6 vssa1
port 643 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 117504 6 vdda2
port 644 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 117504 6 vdda2
port 645 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 117504 6 vdda2
port 646 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 117504 6 vdda2
port 647 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 117504 6 vdda2
port 648 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 117504 6 vdda2
port 649 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 117504 6 vssa2
port 650 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 117504 6 vssa2
port 651 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 117504 6 vssa2
port 652 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 117504 6 vssa2
port 653 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 117504 6 vssa2
port 654 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 117504 6 vssa2
port 655 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 7198572
string GDS_START 339680
<< end >>

